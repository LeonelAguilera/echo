LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY Reg_addr IS
   PORT( 
      sig0 : OUT    std_logic
   );

-- Declarations

END Reg_addr ;

ARCHITECTURE Reg_map OF Reg_addr IS
    
    --signal SDA_data : std_logic_vector
    
BEGIN
END ARCHITECTURE Reg_map;

