--
-- VHDL Architecture echo_lib.parameter_gen.behav
--
-- Created:
--          by - antmo328.student-liu.se (muxen2-112.ad.liu.se)
--          at - 23:11:18 10/12/25
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY parameter_gen IS
-- Declarations

END parameter_gen ;

--
ARCHITECTURE behav OF parameter_gen IS
BEGIN
END ARCHITECTURE behav;

