LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY i2c IS
   PORT( 
      FPGA_clk : IN     std_logic;
      SDA      : OUT    std_logic;
      OK       : OUT    std_logic;
      SCL      : OUT    std_logic;
      Reset    : IN     std_logic;
      Mode     : OUT    std_logic;
      CSB      : OUT    std_logic
   );

-- Declarations

END i2c ;


--
-- VHDL Architecture echo_lib.i2c.struct
--
-- Created:
--          by - alfth698.student-liu.se (muxen2-108.ad.liu.se)
--          at - 14:07:29 10/13/25
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

LIBRARY echo_lib;

ARCHITECTURE struct OF i2c IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL sig0 : std_logic;
   SIGNAL CLK  : std_logic;


   -- Component Declarations
   COMPONENT Clock_div
   PORT (
      FPGA_clk : IN     std_logic ;
      CLK      : OUT    std_logic ;
      Reset    : IN     std_logic 
   );
   END COMPONENT;
   COMPONENT FSM
   PORT (
      Reset : IN     std_logic ;
      sig0  : IN     std_logic 
   );
   END COMPONENT;
   COMPONENT Mode
   PORT (
      Mode : OUT    std_logic ;
      CSB  : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Reg_addr
   PORT (
      sig0 : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT i2c_init
   PORT (
      Reset : IN     std_logic ;
      CLK   : IN     std_logic ;
      SDA   : OUT    std_logic ;
      SCL   : OUT    std_logic ;
      OK    : OUT    std_logic 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Clock_div USE ENTITY echo_lib.Clock_div;
   FOR ALL : FSM USE ENTITY echo_lib.FSM;
   FOR ALL : Mode USE ENTITY echo_lib.Mode;
   FOR ALL : Reg_addr USE ENTITY echo_lib.Reg_addr;
   FOR ALL : i2c_init USE ENTITY echo_lib.i2c_init;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   U_1 : Clock_div
      PORT MAP (
         FPGA_clk => FPGA_clk,
         CLK      => CLK,
         Reset    => Reset
      );
   U_2 : FSM
      PORT MAP (
         Reset => Reset,
         sig0  => sig0
      );
   U_3 : Mode
      PORT MAP (
         Mode => Mode,
         CSB  => CSB
      );
   U_0 : Reg_addr
      PORT MAP (
         sig0 => sig0
      );
   U_4 : i2c_init
      PORT MAP (
         Reset => Reset,
         CLK   => CLK,
         SDA   => SDA,
         SCL   => SCL,
         OK    => OK
      );

END struct;
