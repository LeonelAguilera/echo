--
-- VHDL Architecture echo_lib.i2c.sdfsd
--
-- Created:
--          by - alfth698.student-liu.se (muxen2-116.ad.liu.se)
--          at - 14:21:05 10/16/25
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY i2c IS
   PORT( 
      SDA   : OUT    std_logic;
      SCL   : OUT    std_logic;
      Reset : IN     std_logic;
      HEX6  : OUT    std_logic_vector (0 TO 6);
      HEX7  : OUT    std_logic_vector (0 TO 6);
      c0    : IN     std_logic
   );

-- Declarations

type exemplar_string_array is array (natural range <>, natural range <>) of character;
attribute pin_number : string;
attribute array_pin_number : exemplar_string_array;
attribute array_pin_number of hex6 : signal is ("AC17","AA15","AB15","AB17","AA16","AB16","AA17");
attribute array_pin_number of hex7 : signal is ("AA14","AG18","AF17","AH17","AG17","AE17","AD17");
attribute pin_number of SDA: signal is "A8";
attribute pin_number of SCL: signal is "B7";
attribute pin_number of Reset: signal is "AE14";

END i2c ;

--
-- VHDL Architecture echo_lib.i2c.struct
--
-- Created:
--          by - alfth698.student-liu.se (muxen2-116.ad.liu.se)
--          at - 18:49:48 10/29/25
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

LIBRARY echo_lib;

ARCHITECTURE struct OF i2c IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL CLK_100k : std_logic;
   SIGNAL CLK_200k : std_logic;


   -- Component Declarations
   COMPONENT Clock_div
   PORT (
      CLK_200k : OUT    std_logic ;
      Reset    : IN     std_logic ;
      c0       : IN     std_logic ;
      CLK_100k : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Grp_Nr
   PORT (
      HEX7 : OUT    std_logic_vector (0 TO 6);
      HEX6 : OUT    std_logic_vector (0 TO 6)
   );
   END COMPONENT;
   COMPONENT i2c_init
   PORT (
      Reset    : IN     std_logic ;
      SDA      : OUT    std_logic ;
      SCL      : OUT    std_logic ;
      CLK_200k : IN     std_logic ;
      CLK_100k : IN     std_logic 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Clock_div USE ENTITY echo_lib.Clock_div;
   FOR ALL : Grp_Nr USE ENTITY echo_lib.Grp_Nr;
   FOR ALL : i2c_init USE ENTITY echo_lib.i2c_init;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   U_1 : Clock_div
      PORT MAP (
         CLK_200k => CLK_200k,
         Reset    => Reset,
         c0       => c0,
         CLK_100k => CLK_100k
      );
   U_0 : Grp_Nr
      PORT MAP (
         HEX7 => HEX7,
         HEX6 => HEX6
      );
   U_4 : i2c_init
      PORT MAP (
         Reset    => Reset,
         SDA      => SDA,
         SCL      => SCL,
         CLK_200k => CLK_200k,
         CLK_100k => CLK_100k
      );

END struct;
