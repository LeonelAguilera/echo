LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY i2c IS
   PORT( 
      PLL   : IN     std_logic;
      SDA   : OUT    std_logic;
      SCL   : OUT    std_logic;
      Reset : IN     std_logic
   );

-- Declarations

END i2c ;


--
-- VHDL Architecture echo_lib.i2c.struct
--
-- Created:
--          by - alfth698.student-liu.se (muxen2-116.ad.liu.se)
--          at - 14:48:17 10/16/25
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

LIBRARY echo_lib;

ARCHITECTURE struct OF i2c IS

   -- Architecture declarations
   attribute pin_number of SDA: signal is "A8  ";
   attribute pin_number of SCL: signal is "B7  ";
   attribute pin_number of Reset: signal is "AE14";
   attribute pin_number of PLL : signal is "AF14";

   -- Internal signal declarations
   SIGNAL CLK : std_logic;


type exemplar_string_array is array (natural range <>, natural range <>) of character;
attribute pin_number of SDA: signal is "A8  ";
attribute pin_number of SCL: signal is "B7  ";
attribute pin_number of Reset: signal is "AE14";
attribute pin_number of PLL : signal is "AF14";

   -- Component Declarations
   COMPONENT Clock_div
   PORT (
      CLK   : OUT    std_logic ;
      Reset : IN     std_logic ;
      PLL   : IN     std_logic 
   );
   END COMPONENT;
   COMPONENT i2c_init
   PORT (
      Reset : IN     std_logic ;
      CLK   : IN     std_logic ;
      SDA   : OUT    std_logic ;
      SCL   : OUT    std_logic 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Clock_div USE ENTITY echo_lib.Clock_div;
   FOR ALL : i2c_init USE ENTITY echo_lib.i2c_init;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   U_1 : Clock_div
      PORT MAP (
         CLK   => CLK,
         Reset => Reset,
         PLL   => PLL
      );
   U_4 : i2c_init
      PORT MAP (
         Reset => Reset,
         CLK   => CLK,
         SDA   => SDA,
         SCL   => SCL
      );

END struct;
